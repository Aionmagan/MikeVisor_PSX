pBAV        n      @       �@            �@            �@            �@            �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             @@        ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��               @@        ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��              @@        ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��              @@        ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��              @@        ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��               @@         ��              �?����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    